`timescale 1ns/1ns

module statusRegister (
    input clk, rst,

    input [3:0] status_bits_in,
    input s,
    output reg [3:0] status_bits_out
);

    always @(negedge clk, posedge rst) begin
        if(rst) status_bits_out <= 0;
        else if(s) begin 
            status_bits_out <= status_bits_in;
            $display("%d%d%d%d", status_bits_in[3],status_bits_in[2],status_bits_in[1],status_bits_in[0]);
        end
    end
    
endmodule